`timescale 1ns / 1ps
module i_mem(input [7:0]address, output[31:0]data);
wire [31:0] program[255:0];
assign program[0]=32'b00000000001101101110010000000001;
assign program[1]=32'b00000000001101101110000000011000;
assign program[2]=32'b00000000000100001110000011111111;
assign program[3]=32'b00000010001100001110011100000010;
assign program[4]=32'b00000000001101101110010000000010;
assign program[5]=32'b00000000000001011110000000000001;
assign program[6]=32'b00000001001100001110011100000101;
assign program[7]=32'b00000000001101101110010000000100;
assign program[8]=32'b00000000001101101110000000011000;
assign program[9]=32'b00000000000100001110000011111111;
assign program[10]=32'b00000010001100001110011100001001;
assign program[11]=32'b00000000001101101110010000001000;
assign program[12]=32'b00000000000001011110000000000010;
assign program[13]=32'b00000001001100001110011100001100;
assign program[14]=32'b00000011001101101110011100000000;
assign data=program[address];
endmodule
